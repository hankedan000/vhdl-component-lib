--------------------------------------------------------------------------------
-- Written By: E. George Walters
-- Date Created: 23 Sep 12
-- Last Revision: 23 Sep 12
-- 
-- Entity: BCDAddSUBSlice_tb
-- Description: VHDL test bench for BCDAddSUBSlice.
--
-- Dependencies:
--    BCDAddSubSlice
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.ALL; 
library djh5533_reb5427_Library;
use djh5533_reb5427_Library.djh5533_reb5427_Components.ALL;

--------------------------------------------------------------------------------
entity BCDAddSubSlice_tb is
end BCDAddSubSlice_tb;
--------------------------------------------------------------------------------
 
architecture testbench of BCDAddSubSlice_tb is 
    
   signal A : std_logic_vector(3 downto 0) := (others => '0');
   signal B : std_logic_vector(3 downto 0) := (others => '0');
   signal CBI : std_logic := '0';
   signal SUB : std_logic := '0';

   signal CBO : std_logic;
   signal SUM : std_logic_vector(3 downto 0);
   
   -- Test vector includes input stimuli and expected outputs
   -- A   : bits 14..11
   -- B   : bits 10..7
   -- CBI : bit 6
   -- SUB : bit 5
   -- CBO : bit 4
   -- SUM : bits 3..0
   type test_vector_type is array (0 to 399) of std_logic_vector(14 downto 0); -- test vector is A & B & CBI & SUM & CBO & SUM
   constant test_vector : test_vector_type := (
      -- A        B     CBI   SUB   CBO    SUM
      "0000" & "0000" & '0' & '0' & '0' & "0000",
      "0000" & "0001" & '0' & '0' & '0' & "0001",
      "0000" & "0010" & '0' & '0' & '0' & "0010",
      "0000" & "0011" & '0' & '0' & '0' & "0011",
      "0000" & "0100" & '0' & '0' & '0' & "0100",
      "0000" & "0101" & '0' & '0' & '0' & "0101",
      "0000" & "0110" & '0' & '0' & '0' & "0110",
      "0000" & "0111" & '0' & '0' & '0' & "0111",
      "0000" & "1000" & '0' & '0' & '0' & "1000",
      "0000" & "1001" & '0' & '0' & '0' & "1001",
      "0001" & "0000" & '0' & '0' & '0' & "0001",
      "0001" & "0001" & '0' & '0' & '0' & "0010",
      "0001" & "0010" & '0' & '0' & '0' & "0011",
      "0001" & "0011" & '0' & '0' & '0' & "0100",
      "0001" & "0100" & '0' & '0' & '0' & "0101",
      "0001" & "0101" & '0' & '0' & '0' & "0110",
      "0001" & "0110" & '0' & '0' & '0' & "0111",
      "0001" & "0111" & '0' & '0' & '0' & "1000",
      "0001" & "1000" & '0' & '0' & '0' & "1001",
      "0001" & "1001" & '0' & '0' & '1' & "0000",
      "0010" & "0000" & '0' & '0' & '0' & "0010",
      "0010" & "0001" & '0' & '0' & '0' & "0011",
      "0010" & "0010" & '0' & '0' & '0' & "0100",
      "0010" & "0011" & '0' & '0' & '0' & "0101",
      "0010" & "0100" & '0' & '0' & '0' & "0110",
      "0010" & "0101" & '0' & '0' & '0' & "0111",
      "0010" & "0110" & '0' & '0' & '0' & "1000",
      "0010" & "0111" & '0' & '0' & '0' & "1001",
      "0010" & "1000" & '0' & '0' & '1' & "0000",
      "0010" & "1001" & '0' & '0' & '1' & "0001",
      "0011" & "0000" & '0' & '0' & '0' & "0011",
      "0011" & "0001" & '0' & '0' & '0' & "0100",
      "0011" & "0010" & '0' & '0' & '0' & "0101",
      "0011" & "0011" & '0' & '0' & '0' & "0110",
      "0011" & "0100" & '0' & '0' & '0' & "0111",
      "0011" & "0101" & '0' & '0' & '0' & "1000",
      "0011" & "0110" & '0' & '0' & '0' & "1001",
      "0011" & "0111" & '0' & '0' & '1' & "0000",
      "0011" & "1000" & '0' & '0' & '1' & "0001",
      "0011" & "1001" & '0' & '0' & '1' & "0010",
      "0100" & "0000" & '0' & '0' & '0' & "0100",
      "0100" & "0001" & '0' & '0' & '0' & "0101",
      "0100" & "0010" & '0' & '0' & '0' & "0110",
      "0100" & "0011" & '0' & '0' & '0' & "0111",
      "0100" & "0100" & '0' & '0' & '0' & "1000",
      "0100" & "0101" & '0' & '0' & '0' & "1001",
      "0100" & "0110" & '0' & '0' & '1' & "0000",
      "0100" & "0111" & '0' & '0' & '1' & "0001",
      "0100" & "1000" & '0' & '0' & '1' & "0010",
      "0100" & "1001" & '0' & '0' & '1' & "0011",
      "0101" & "0000" & '0' & '0' & '0' & "0101",
      "0101" & "0001" & '0' & '0' & '0' & "0110",
      "0101" & "0010" & '0' & '0' & '0' & "0111",
      "0101" & "0011" & '0' & '0' & '0' & "1000",
      "0101" & "0100" & '0' & '0' & '0' & "1001",
      "0101" & "0101" & '0' & '0' & '1' & "0000",
      "0101" & "0110" & '0' & '0' & '1' & "0001",
      "0101" & "0111" & '0' & '0' & '1' & "0010",
      "0101" & "1000" & '0' & '0' & '1' & "0011",
      "0101" & "1001" & '0' & '0' & '1' & "0100",
      "0110" & "0000" & '0' & '0' & '0' & "0110",
      "0110" & "0001" & '0' & '0' & '0' & "0111",
      "0110" & "0010" & '0' & '0' & '0' & "1000",
      "0110" & "0011" & '0' & '0' & '0' & "1001",
      "0110" & "0100" & '0' & '0' & '1' & "0000",
      "0110" & "0101" & '0' & '0' & '1' & "0001",
      "0110" & "0110" & '0' & '0' & '1' & "0010",
      "0110" & "0111" & '0' & '0' & '1' & "0011",
      "0110" & "1000" & '0' & '0' & '1' & "0100",
      "0110" & "1001" & '0' & '0' & '1' & "0101",
      "0111" & "0000" & '0' & '0' & '0' & "0111",
      "0111" & "0001" & '0' & '0' & '0' & "1000",
      "0111" & "0010" & '0' & '0' & '0' & "1001",
      "0111" & "0011" & '0' & '0' & '1' & "0000",
      "0111" & "0100" & '0' & '0' & '1' & "0001",
      "0111" & "0101" & '0' & '0' & '1' & "0010",
      "0111" & "0110" & '0' & '0' & '1' & "0011",
      "0111" & "0111" & '0' & '0' & '1' & "0100",
      "0111" & "1000" & '0' & '0' & '1' & "0101",
      "0111" & "1001" & '0' & '0' & '1' & "0110",
      "1000" & "0000" & '0' & '0' & '0' & "1000",
      "1000" & "0001" & '0' & '0' & '0' & "1001",
      "1000" & "0010" & '0' & '0' & '1' & "0000",
      "1000" & "0011" & '0' & '0' & '1' & "0001",
      "1000" & "0100" & '0' & '0' & '1' & "0010",
      "1000" & "0101" & '0' & '0' & '1' & "0011",
      "1000" & "0110" & '0' & '0' & '1' & "0100",
      "1000" & "0111" & '0' & '0' & '1' & "0101",
      "1000" & "1000" & '0' & '0' & '1' & "0110",
      "1000" & "1001" & '0' & '0' & '1' & "0111",
      "1001" & "0000" & '0' & '0' & '0' & "1001",
      "1001" & "0001" & '0' & '0' & '1' & "0000",
      "1001" & "0010" & '0' & '0' & '1' & "0001",
      "1001" & "0011" & '0' & '0' & '1' & "0010",
      "1001" & "0100" & '0' & '0' & '1' & "0011",
      "1001" & "0101" & '0' & '0' & '1' & "0100",
      "1001" & "0110" & '0' & '0' & '1' & "0101",
      "1001" & "0111" & '0' & '0' & '1' & "0110",
      "1001" & "1000" & '0' & '0' & '1' & "0111",
      "1001" & "1001" & '0' & '0' & '1' & "1000",
      "0000" & "0000" & '0' & '1' & '0' & "0000",
      "0000" & "0001" & '0' & '1' & '1' & "1001",
      "0000" & "0010" & '0' & '1' & '1' & "1000",
      "0000" & "0011" & '0' & '1' & '1' & "0111",
      "0000" & "0100" & '0' & '1' & '1' & "0110",
      "0000" & "0101" & '0' & '1' & '1' & "0101",
      "0000" & "0110" & '0' & '1' & '1' & "0100",
      "0000" & "0111" & '0' & '1' & '1' & "0011",
      "0000" & "1000" & '0' & '1' & '1' & "0010",
      "0000" & "1001" & '0' & '1' & '1' & "0001",
      "0001" & "0000" & '0' & '1' & '0' & "0001",
      "0001" & "0001" & '0' & '1' & '0' & "0000",
      "0001" & "0010" & '0' & '1' & '1' & "1001",
      "0001" & "0011" & '0' & '1' & '1' & "1000",
      "0001" & "0100" & '0' & '1' & '1' & "0111",
      "0001" & "0101" & '0' & '1' & '1' & "0110",
      "0001" & "0110" & '0' & '1' & '1' & "0101",
      "0001" & "0111" & '0' & '1' & '1' & "0100",
      "0001" & "1000" & '0' & '1' & '1' & "0011",
      "0001" & "1001" & '0' & '1' & '1' & "0010",
      "0010" & "0000" & '0' & '1' & '0' & "0010",
      "0010" & "0001" & '0' & '1' & '0' & "0001",
      "0010" & "0010" & '0' & '1' & '0' & "0000",
      "0010" & "0011" & '0' & '1' & '1' & "1001",
      "0010" & "0100" & '0' & '1' & '1' & "1000",
      "0010" & "0101" & '0' & '1' & '1' & "0111",
      "0010" & "0110" & '0' & '1' & '1' & "0110",
      "0010" & "0111" & '0' & '1' & '1' & "0101",
      "0010" & "1000" & '0' & '1' & '1' & "0100",
      "0010" & "1001" & '0' & '1' & '1' & "0011",
      "0011" & "0000" & '0' & '1' & '0' & "0011",
      "0011" & "0001" & '0' & '1' & '0' & "0010",
      "0011" & "0010" & '0' & '1' & '0' & "0001",
      "0011" & "0011" & '0' & '1' & '0' & "0000",
      "0011" & "0100" & '0' & '1' & '1' & "1001",
      "0011" & "0101" & '0' & '1' & '1' & "1000",
      "0011" & "0110" & '0' & '1' & '1' & "0111",
      "0011" & "0111" & '0' & '1' & '1' & "0110",
      "0011" & "1000" & '0' & '1' & '1' & "0101",
      "0011" & "1001" & '0' & '1' & '1' & "0100",
      "0100" & "0000" & '0' & '1' & '0' & "0100",
      "0100" & "0001" & '0' & '1' & '0' & "0011",
      "0100" & "0010" & '0' & '1' & '0' & "0010",
      "0100" & "0011" & '0' & '1' & '0' & "0001",
      "0100" & "0100" & '0' & '1' & '0' & "0000",
      "0100" & "0101" & '0' & '1' & '1' & "1001",
      "0100" & "0110" & '0' & '1' & '1' & "1000",
      "0100" & "0111" & '0' & '1' & '1' & "0111",
      "0100" & "1000" & '0' & '1' & '1' & "0110",
      "0100" & "1001" & '0' & '1' & '1' & "0101",
      "0101" & "0000" & '0' & '1' & '0' & "0101",
      "0101" & "0001" & '0' & '1' & '0' & "0100",
      "0101" & "0010" & '0' & '1' & '0' & "0011",
      "0101" & "0011" & '0' & '1' & '0' & "0010",
      "0101" & "0100" & '0' & '1' & '0' & "0001",
      "0101" & "0101" & '0' & '1' & '0' & "0000",
      "0101" & "0110" & '0' & '1' & '1' & "1001",
      "0101" & "0111" & '0' & '1' & '1' & "1000",
      "0101" & "1000" & '0' & '1' & '1' & "0111",
      "0101" & "1001" & '0' & '1' & '1' & "0110",
      "0110" & "0000" & '0' & '1' & '0' & "0110",
      "0110" & "0001" & '0' & '1' & '0' & "0101",
      "0110" & "0010" & '0' & '1' & '0' & "0100",
      "0110" & "0011" & '0' & '1' & '0' & "0011",
      "0110" & "0100" & '0' & '1' & '0' & "0010",
      "0110" & "0101" & '0' & '1' & '0' & "0001",
      "0110" & "0110" & '0' & '1' & '0' & "0000",
      "0110" & "0111" & '0' & '1' & '1' & "1001",
      "0110" & "1000" & '0' & '1' & '1' & "1000",
      "0110" & "1001" & '0' & '1' & '1' & "0111",
      "0111" & "0000" & '0' & '1' & '0' & "0111",
      "0111" & "0001" & '0' & '1' & '0' & "0110",
      "0111" & "0010" & '0' & '1' & '0' & "0101",
      "0111" & "0011" & '0' & '1' & '0' & "0100",
      "0111" & "0100" & '0' & '1' & '0' & "0011",
      "0111" & "0101" & '0' & '1' & '0' & "0010",
      "0111" & "0110" & '0' & '1' & '0' & "0001",
      "0111" & "0111" & '0' & '1' & '0' & "0000",
      "0111" & "1000" & '0' & '1' & '1' & "1001",
      "0111" & "1001" & '0' & '1' & '1' & "1000",
      "1000" & "0000" & '0' & '1' & '0' & "1000",
      "1000" & "0001" & '0' & '1' & '0' & "0111",
      "1000" & "0010" & '0' & '1' & '0' & "0110",
      "1000" & "0011" & '0' & '1' & '0' & "0101",
      "1000" & "0100" & '0' & '1' & '0' & "0100",
      "1000" & "0101" & '0' & '1' & '0' & "0011",
      "1000" & "0110" & '0' & '1' & '0' & "0010",
      "1000" & "0111" & '0' & '1' & '0' & "0001",
      "1000" & "1000" & '0' & '1' & '0' & "0000",
      "1000" & "1001" & '0' & '1' & '1' & "1001",
      "1001" & "0000" & '0' & '1' & '0' & "1001",
      "1001" & "0001" & '0' & '1' & '0' & "1000",
      "1001" & "0010" & '0' & '1' & '0' & "0111",
      "1001" & "0011" & '0' & '1' & '0' & "0110",
      "1001" & "0100" & '0' & '1' & '0' & "0101",
      "1001" & "0101" & '0' & '1' & '0' & "0100",
      "1001" & "0110" & '0' & '1' & '0' & "0011",
      "1001" & "0111" & '0' & '1' & '0' & "0010",
      "1001" & "1000" & '0' & '1' & '0' & "0001",
      "1001" & "1001" & '0' & '1' & '0' & "0000",
      "0000" & "0000" & '1' & '0' & '0' & "0001",
      "0000" & "0001" & '1' & '0' & '0' & "0010",
      "0000" & "0010" & '1' & '0' & '0' & "0011",
      "0000" & "0011" & '1' & '0' & '0' & "0100",
      "0000" & "0100" & '1' & '0' & '0' & "0101",
      "0000" & "0101" & '1' & '0' & '0' & "0110",
      "0000" & "0110" & '1' & '0' & '0' & "0111",
      "0000" & "0111" & '1' & '0' & '0' & "1000",
      "0000" & "1000" & '1' & '0' & '0' & "1001",
      "0000" & "1001" & '1' & '0' & '1' & "0000",
      "0001" & "0000" & '1' & '0' & '0' & "0010",
      "0001" & "0001" & '1' & '0' & '0' & "0011",
      "0001" & "0010" & '1' & '0' & '0' & "0100",
      "0001" & "0011" & '1' & '0' & '0' & "0101",
      "0001" & "0100" & '1' & '0' & '0' & "0110",
      "0001" & "0101" & '1' & '0' & '0' & "0111",
      "0001" & "0110" & '1' & '0' & '0' & "1000",
      "0001" & "0111" & '1' & '0' & '0' & "1001",
      "0001" & "1000" & '1' & '0' & '1' & "0000",
      "0001" & "1001" & '1' & '0' & '1' & "0001",
      "0010" & "0000" & '1' & '0' & '0' & "0011",
      "0010" & "0001" & '1' & '0' & '0' & "0100",
      "0010" & "0010" & '1' & '0' & '0' & "0101",
      "0010" & "0011" & '1' & '0' & '0' & "0110",
      "0010" & "0100" & '1' & '0' & '0' & "0111",
      "0010" & "0101" & '1' & '0' & '0' & "1000",
      "0010" & "0110" & '1' & '0' & '0' & "1001",
      "0010" & "0111" & '1' & '0' & '1' & "0000",
      "0010" & "1000" & '1' & '0' & '1' & "0001",
      "0010" & "1001" & '1' & '0' & '1' & "0010",
      "0011" & "0000" & '1' & '0' & '0' & "0100",
      "0011" & "0001" & '1' & '0' & '0' & "0101",
      "0011" & "0010" & '1' & '0' & '0' & "0110",
      "0011" & "0011" & '1' & '0' & '0' & "0111",
      "0011" & "0100" & '1' & '0' & '0' & "1000",
      "0011" & "0101" & '1' & '0' & '0' & "1001",
      "0011" & "0110" & '1' & '0' & '1' & "0000",
      "0011" & "0111" & '1' & '0' & '1' & "0001",
      "0011" & "1000" & '1' & '0' & '1' & "0010",
      "0011" & "1001" & '1' & '0' & '1' & "0011",
      "0100" & "0000" & '1' & '0' & '0' & "0101",
      "0100" & "0001" & '1' & '0' & '0' & "0110",
      "0100" & "0010" & '1' & '0' & '0' & "0111",
      "0100" & "0011" & '1' & '0' & '0' & "1000",
      "0100" & "0100" & '1' & '0' & '0' & "1001",
      "0100" & "0101" & '1' & '0' & '1' & "0000",
      "0100" & "0110" & '1' & '0' & '1' & "0001",
      "0100" & "0111" & '1' & '0' & '1' & "0010",
      "0100" & "1000" & '1' & '0' & '1' & "0011",
      "0100" & "1001" & '1' & '0' & '1' & "0100",
      "0101" & "0000" & '1' & '0' & '0' & "0110",
      "0101" & "0001" & '1' & '0' & '0' & "0111",
      "0101" & "0010" & '1' & '0' & '0' & "1000",
      "0101" & "0011" & '1' & '0' & '0' & "1001",
      "0101" & "0100" & '1' & '0' & '1' & "0000",
      "0101" & "0101" & '1' & '0' & '1' & "0001",
      "0101" & "0110" & '1' & '0' & '1' & "0010",
      "0101" & "0111" & '1' & '0' & '1' & "0011",
      "0101" & "1000" & '1' & '0' & '1' & "0100",
      "0101" & "1001" & '1' & '0' & '1' & "0101",
      "0110" & "0000" & '1' & '0' & '0' & "0111",
      "0110" & "0001" & '1' & '0' & '0' & "1000",
      "0110" & "0010" & '1' & '0' & '0' & "1001",
      "0110" & "0011" & '1' & '0' & '1' & "0000",
      "0110" & "0100" & '1' & '0' & '1' & "0001",
      "0110" & "0101" & '1' & '0' & '1' & "0010",
      "0110" & "0110" & '1' & '0' & '1' & "0011",
      "0110" & "0111" & '1' & '0' & '1' & "0100",
      "0110" & "1000" & '1' & '0' & '1' & "0101",
      "0110" & "1001" & '1' & '0' & '1' & "0110",
      "0111" & "0000" & '1' & '0' & '0' & "1000",
      "0111" & "0001" & '1' & '0' & '0' & "1001",
      "0111" & "0010" & '1' & '0' & '1' & "0000",
      "0111" & "0011" & '1' & '0' & '1' & "0001",
      "0111" & "0100" & '1' & '0' & '1' & "0010",
      "0111" & "0101" & '1' & '0' & '1' & "0011",
      "0111" & "0110" & '1' & '0' & '1' & "0100",
      "0111" & "0111" & '1' & '0' & '1' & "0101",
      "0111" & "1000" & '1' & '0' & '1' & "0110",
      "0111" & "1001" & '1' & '0' & '1' & "0111",
      "1000" & "0000" & '1' & '0' & '0' & "1001",
      "1000" & "0001" & '1' & '0' & '1' & "0000",
      "1000" & "0010" & '1' & '0' & '1' & "0001",
      "1000" & "0011" & '1' & '0' & '1' & "0010",
      "1000" & "0100" & '1' & '0' & '1' & "0011",
      "1000" & "0101" & '1' & '0' & '1' & "0100",
      "1000" & "0110" & '1' & '0' & '1' & "0101",
      "1000" & "0111" & '1' & '0' & '1' & "0110",
      "1000" & "1000" & '1' & '0' & '1' & "0111",
      "1000" & "1001" & '1' & '0' & '1' & "1000",
      "1001" & "0000" & '1' & '0' & '1' & "0000",
      "1001" & "0001" & '1' & '0' & '1' & "0001",
      "1001" & "0010" & '1' & '0' & '1' & "0010",
      "1001" & "0011" & '1' & '0' & '1' & "0011",
      "1001" & "0100" & '1' & '0' & '1' & "0100",
      "1001" & "0101" & '1' & '0' & '1' & "0101",
      "1001" & "0110" & '1' & '0' & '1' & "0110",
      "1001" & "0111" & '1' & '0' & '1' & "0111",
      "1001" & "1000" & '1' & '0' & '1' & "1000",
      "1001" & "1001" & '1' & '0' & '1' & "1001",
      "0000" & "0000" & '1' & '1' & '1' & "1001",
      "0000" & "0001" & '1' & '1' & '1' & "1000",
      "0000" & "0010" & '1' & '1' & '1' & "0111",
      "0000" & "0011" & '1' & '1' & '1' & "0110",
      "0000" & "0100" & '1' & '1' & '1' & "0101",
      "0000" & "0101" & '1' & '1' & '1' & "0100",
      "0000" & "0110" & '1' & '1' & '1' & "0011",
      "0000" & "0111" & '1' & '1' & '1' & "0010",
      "0000" & "1000" & '1' & '1' & '1' & "0001",
      "0000" & "1001" & '1' & '1' & '1' & "0000",
      "0001" & "0000" & '1' & '1' & '0' & "0000",
      "0001" & "0001" & '1' & '1' & '1' & "1001",
      "0001" & "0010" & '1' & '1' & '1' & "1000",
      "0001" & "0011" & '1' & '1' & '1' & "0111",
      "0001" & "0100" & '1' & '1' & '1' & "0110",
      "0001" & "0101" & '1' & '1' & '1' & "0101",
      "0001" & "0110" & '1' & '1' & '1' & "0100",
      "0001" & "0111" & '1' & '1' & '1' & "0011",
      "0001" & "1000" & '1' & '1' & '1' & "0010",
      "0001" & "1001" & '1' & '1' & '1' & "0001",
      "0010" & "0000" & '1' & '1' & '0' & "0001",
      "0010" & "0001" & '1' & '1' & '0' & "0000",
      "0010" & "0010" & '1' & '1' & '1' & "1001",
      "0010" & "0011" & '1' & '1' & '1' & "1000",
      "0010" & "0100" & '1' & '1' & '1' & "0111",
      "0010" & "0101" & '1' & '1' & '1' & "0110",
      "0010" & "0110" & '1' & '1' & '1' & "0101",
      "0010" & "0111" & '1' & '1' & '1' & "0100",
      "0010" & "1000" & '1' & '1' & '1' & "0011",
      "0010" & "1001" & '1' & '1' & '1' & "0010",
      "0011" & "0000" & '1' & '1' & '0' & "0010",
      "0011" & "0001" & '1' & '1' & '0' & "0001",
      "0011" & "0010" & '1' & '1' & '0' & "0000",
      "0011" & "0011" & '1' & '1' & '1' & "1001",
      "0011" & "0100" & '1' & '1' & '1' & "1000",
      "0011" & "0101" & '1' & '1' & '1' & "0111",
      "0011" & "0110" & '1' & '1' & '1' & "0110",
      "0011" & "0111" & '1' & '1' & '1' & "0101",
      "0011" & "1000" & '1' & '1' & '1' & "0100",
      "0011" & "1001" & '1' & '1' & '1' & "0011",
      "0100" & "0000" & '1' & '1' & '0' & "0011",
      "0100" & "0001" & '1' & '1' & '0' & "0010",
      "0100" & "0010" & '1' & '1' & '0' & "0001",
      "0100" & "0011" & '1' & '1' & '0' & "0000",
      "0100" & "0100" & '1' & '1' & '1' & "1001",
      "0100" & "0101" & '1' & '1' & '1' & "1000",
      "0100" & "0110" & '1' & '1' & '1' & "0111",
      "0100" & "0111" & '1' & '1' & '1' & "0110",
      "0100" & "1000" & '1' & '1' & '1' & "0101",
      "0100" & "1001" & '1' & '1' & '1' & "0100",
      "0101" & "0000" & '1' & '1' & '0' & "0100",
      "0101" & "0001" & '1' & '1' & '0' & "0011",
      "0101" & "0010" & '1' & '1' & '0' & "0010",
      "0101" & "0011" & '1' & '1' & '0' & "0001",
      "0101" & "0100" & '1' & '1' & '0' & "0000",
      "0101" & "0101" & '1' & '1' & '1' & "1001",
      "0101" & "0110" & '1' & '1' & '1' & "1000",
      "0101" & "0111" & '1' & '1' & '1' & "0111",
      "0101" & "1000" & '1' & '1' & '1' & "0110",
      "0101" & "1001" & '1' & '1' & '1' & "0101",
      "0110" & "0000" & '1' & '1' & '0' & "0101",
      "0110" & "0001" & '1' & '1' & '0' & "0100",
      "0110" & "0010" & '1' & '1' & '0' & "0011",
      "0110" & "0011" & '1' & '1' & '0' & "0010",
      "0110" & "0100" & '1' & '1' & '0' & "0001",
      "0110" & "0101" & '1' & '1' & '0' & "0000",
      "0110" & "0110" & '1' & '1' & '1' & "1001",
      "0110" & "0111" & '1' & '1' & '1' & "1000",
      "0110" & "1000" & '1' & '1' & '1' & "0111",
      "0110" & "1001" & '1' & '1' & '1' & "0110",
      "0111" & "0000" & '1' & '1' & '0' & "0110",
      "0111" & "0001" & '1' & '1' & '0' & "0101",
      "0111" & "0010" & '1' & '1' & '0' & "0100",
      "0111" & "0011" & '1' & '1' & '0' & "0011",
      "0111" & "0100" & '1' & '1' & '0' & "0010",
      "0111" & "0101" & '1' & '1' & '0' & "0001",
      "0111" & "0110" & '1' & '1' & '0' & "0000",
      "0111" & "0111" & '1' & '1' & '1' & "1001",
      "0111" & "1000" & '1' & '1' & '1' & "1000",
      "0111" & "1001" & '1' & '1' & '1' & "0111",
      "1000" & "0000" & '1' & '1' & '0' & "0111",
      "1000" & "0001" & '1' & '1' & '0' & "0110",
      "1000" & "0010" & '1' & '1' & '0' & "0101",
      "1000" & "0011" & '1' & '1' & '0' & "0100",
      "1000" & "0100" & '1' & '1' & '0' & "0011",
      "1000" & "0101" & '1' & '1' & '0' & "0010",
      "1000" & "0110" & '1' & '1' & '0' & "0001",
      "1000" & "0111" & '1' & '1' & '0' & "0000",
      "1000" & "1000" & '1' & '1' & '1' & "1001",
      "1000" & "1001" & '1' & '1' & '1' & "1000",
      "1001" & "0000" & '1' & '1' & '0' & "1000",
      "1001" & "0001" & '1' & '1' & '0' & "0111",
      "1001" & "0010" & '1' & '1' & '0' & "0110",
      "1001" & "0011" & '1' & '1' & '0' & "0101",
      "1001" & "0100" & '1' & '1' & '0' & "0100",
      "1001" & "0101" & '1' & '1' & '0' & "0011",
      "1001" & "0110" & '1' & '1' & '0' & "0010",
      "1001" & "0111" & '1' & '1' & '0' & "0001",
      "1001" & "1000" & '1' & '1' & '0' & "0000",
      "1001" & "1001" & '1' & '1' & '1' & "1001"
   );
 
begin

   uut: BCDAddSubSlice port map (A, B, CBI, SUB, CBO, SUM);

   process
   begin
      for i in test_vector'Range loop
      
         -- Assign test inputs
         A <= test_vector(i)(14 downto 11);
         B <= test_vector(i)(10 downto 7);
         CBI <= test_vector(i)(6);
         SUB <= test_vector(i)(5);
         
         -- Compare outputs to expected values
         wait for 2ns;
         assert (CBO = test_vector(i)(4) and SUM = test_vector(i)(3 downto 0))
            report "***** Test failed. *****"
            severity Failure;
      end loop;
      
      -- All tests are successful if we get this far
      report "***** All tests completed successfully. *****";
      wait;
   end process;

end testbench;
