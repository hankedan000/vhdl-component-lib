----------------------------------------------------------------------------
-- Entity:        Decoder3to8
-- Written By:    Daniel Hankewycz & Robby Brague
-- Date Created:  9/11/2014
-- Description:   Implements a 3 to 8 bit decoder
--
-- Revision History (date, initials, description):
-- 
-- Dependencies:
--		Mux4to1
----------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity Decoder3to8 is
    Port ( 	X			:	in		STD_LOGIC_VECTOR (2 downto 0);
				EN			:	in		STD_LOGIC;
			  
				Y			: 	out	STD_LOGIC_VECTOR (7 downto 0));
end Decoder3to8;

architecture dataflow of Decoder3to8 is
signal	y_mux	:	STD_LOGIC_VECTOR	(7 downto 0);

begin
	with EN select
		Y	<=	y_mux when '1',
				x"00"	when others;

	with X select
		y_mux <=	"00000001" when "000",
					"00000010" when "001",
					"00000100" when "010",
					"00001000" when "011",
					"00010000" when "100",
					"00100000" when "101",
					"01000000" when "110",
					"10000000" when "111",
					"00000000" when others;
	
end dataflow;