--------------------------------------------------------------------------------
-- Written By: E. George Walters
-- Date Created: 23 Sep 12
-- Last Revision: 23 Sep 12
-- 
-- Entity: BCD_AddSub_tb
-- Description: VHDL test bench for BCD_AddSub.
--
-- Dependencies:
--    BCD_AddSubSlice
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.ALL; 
library djh5533_reb5427_Library;
use djh5533_reb5427_Library.djh5533_reb5427_Components.ALL;

--------------------------------------------------------------------------------
entity BCD_AddSub_tb is
end BCD_AddSub_tb;
--------------------------------------------------------------------------------
 
architecture testbench of BCD_AddSub_tb is 

   signal A : std_logic_vector(15 downto 0) := (others => '0');
   signal B : std_logic_vector(15 downto 0) := (others => '0');
   signal cbi : std_logic := '0';
   signal sub : std_logic := '0';

   signal cbo : std_logic;
   signal sum : std_logic_vector(15 downto 0);
   
   -- Test vector includes input stimuli and expected outputs
   -- A   : bits 50..35
   -- B   : bits 34..19
   -- cbi : bit 18
   -- sub : bit 17
   -- cbo : bit 16
   -- sum : bits 15..0
   type test_vector_type is array (0 to 199) of std_logic_vector(50 downto 0); -- test vector is A & B & cbi & sub & cbo & sum
   constant test_vector : test_vector_type := (
      -- A        B     cbi   sum   cbo    sum
      x"0000" & x"0000" & '0' & '0' & '0' & x"0000",
      x"0000" & x"0001" & '0' & '0' & '0' & x"0001",
      x"0001" & x"0000" & '0' & '0' & '0' & x"0001",
      x"0001" & x"0001" & '0' & '0' & '0' & x"0002",
      x"0009" & x"0001" & '0' & '0' & '0' & x"0010",
      x"9999" & x"0001" & '0' & '0' & '1' & x"0000",
      x"9999" & x"1111" & '0' & '0' & '1' & x"1110",
      x"9000" & x"1000" & '0' & '0' & '1' & x"0000",
      x"0001" & x"0009" & '0' & '0' & '0' & x"0010",
      x"0001" & x"9999" & '0' & '0' & '1' & x"0000",
      x"1111" & x"9999" & '0' & '0' & '1' & x"1110",
      x"1000" & x"9000" & '0' & '0' & '1' & x"0000",
      x"0000" & x"0000" & '0' & '1' & '0' & x"0000",
      x"0000" & x"0001" & '0' & '1' & '1' & x"9999",
      x"0001" & x"0000" & '0' & '1' & '0' & x"0001",
      x"0001" & x"0001" & '0' & '1' & '0' & x"0000",
      x"0009" & x"0001" & '0' & '1' & '0' & x"0008",
      x"9999" & x"0001" & '0' & '1' & '0' & x"9998",
      x"9999" & x"1111" & '0' & '1' & '0' & x"8888",
      x"9000" & x"1000" & '0' & '1' & '0' & x"8000",
      x"0001" & x"0009" & '0' & '1' & '1' & x"9992",
      x"0001" & x"9999" & '0' & '1' & '1' & x"0002",
      x"1111" & x"9999" & '0' & '1' & '1' & x"1112",
      x"1000" & x"9000" & '0' & '1' & '1' & x"2000",
      x"0000" & x"0000" & '1' & '0' & '0' & x"0001",
      x"0000" & x"0001" & '1' & '0' & '0' & x"0002",
      x"0001" & x"0000" & '1' & '0' & '0' & x"0002",
      x"0001" & x"0001" & '1' & '0' & '0' & x"0003",
      x"0009" & x"0001" & '1' & '0' & '0' & x"0011",
      x"9999" & x"0001" & '1' & '0' & '1' & x"0001",
      x"9999" & x"1111" & '1' & '0' & '1' & x"1111",
      x"9000" & x"1000" & '1' & '0' & '1' & x"0001",
      x"0001" & x"0009" & '1' & '0' & '0' & x"0011",
      x"0001" & x"9999" & '1' & '0' & '1' & x"0001",
      x"1111" & x"9999" & '1' & '0' & '1' & x"1111",
      x"1000" & x"9000" & '1' & '0' & '1' & x"0001",
      x"0000" & x"0000" & '1' & '1' & '1' & x"9999",
      x"0000" & x"0001" & '1' & '1' & '1' & x"9998",
      x"0001" & x"0000" & '1' & '1' & '0' & x"0000",
      x"0001" & x"0001" & '1' & '1' & '1' & x"9999",
      x"0009" & x"0001" & '1' & '1' & '0' & x"0007",
      x"9999" & x"0001" & '1' & '1' & '0' & x"9997",
      x"9999" & x"1111" & '1' & '1' & '0' & x"8887",
      x"9000" & x"1000" & '1' & '1' & '0' & x"7999",
      x"0001" & x"0009" & '1' & '1' & '1' & x"9991",
      x"0001" & x"9999" & '1' & '1' & '1' & x"0001",
      x"1111" & x"9999" & '1' & '1' & '1' & x"1111",
      x"1000" & x"9000" & '1' & '1' & '1' & x"1999",
      x"8780" & x"1709" & '0' & '1' & '0' & x"7071",
      x"1125" & x"6327" & '0' & '0' & '0' & x"7452",
      x"0004" & x"6971" & '0' & '1' & '1' & x"3033",
      x"5606" & x"3206" & '0' & '0' & '0' & x"8812",
      x"5794" & x"0087" & '0' & '0' & '0' & x"5881",
      x"9096" & x"5468" & '1' & '0' & '1' & x"4565",
      x"4728" & x"2993" & '0' & '0' & '0' & x"7721",
      x"1376" & x"9851" & '1' & '0' & '1' & x"1228",
      x"5473" & x"6887" & '0' & '0' & '1' & x"2360",
      x"9447" & x"2103" & '1' & '0' & '1' & x"1551",
      x"2547" & x"7057" & '0' & '0' & '0' & x"9604",
      x"9388" & x"2985" & '0' & '1' & '0' & x"6403",
      x"9233" & x"7324" & '0' & '1' & '0' & x"1909",
      x"7637" & x"4069" & '1' & '0' & '1' & x"1707",
      x"3387" & x"9599" & '0' & '0' & '1' & x"2986",
      x"8065" & x"6540" & '0' & '0' & '1' & x"4605",
      x"1191" & x"4477" & '1' & '0' & '0' & x"5669",
      x"6508" & x"7454" & '1' & '0' & '1' & x"3963",
      x"8312" & x"3856" & '1' & '1' & '0' & x"4455",
      x"3018" & x"1882" & '0' & '0' & '0' & x"4900",
      x"2467" & x"8621" & '1' & '1' & '1' & x"3845",
      x"5476" & x"8596" & '0' & '1' & '1' & x"6880",
      x"7580" & x"1302" & '0' & '0' & '0' & x"8882",
      x"8578" & x"1281" & '1' & '0' & '0' & x"9860",
      x"0782" & x"6123" & '0' & '0' & '0' & x"6905",
      x"7259" & x"6512" & '0' & '1' & '0' & x"0747",
      x"4967" & x"1723" & '0' & '0' & '0' & x"6690",
      x"3344" & x"8363" & '0' & '0' & '1' & x"1707",
      x"0583" & x"8527" & '0' & '1' & '1' & x"2056",
      x"8568" & x"2681" & '1' & '0' & '1' & x"1250",
      x"7430" & x"0282" & '1' & '1' & '0' & x"7147",
      x"2397" & x"8527" & '0' & '1' & '1' & x"3870",
      x"0718" & x"9127" & '0' & '1' & '1' & x"1591",
      x"8898" & x"5001" & '0' & '0' & '1' & x"3899",
      x"2256" & x"4843" & '1' & '1' & '1' & x"7412",
      x"0976" & x"0248" & '0' & '0' & '0' & x"1224",
      x"1239" & x"8841" & '1' & '1' & '1' & x"2397",
      x"2208" & x"6687" & '1' & '1' & '1' & x"5520",
      x"4472" & x"8173" & '1' & '1' & '1' & x"6298",
      x"4924" & x"8495" & '1' & '1' & '1' & x"6428",
      x"4281" & x"8021" & '0' & '0' & '1' & x"2302",
      x"1530" & x"3719" & '1' & '1' & '1' & x"7810",
      x"1956" & x"5535" & '0' & '1' & '1' & x"6421",
      x"7449" & x"2689" & '0' & '1' & '0' & x"4760",
      x"6468" & x"6913" & '0' & '1' & '1' & x"9555",
      x"4116" & x"5730" & '0' & '0' & '0' & x"9846",
      x"9716" & x"4392" & '0' & '0' & '1' & x"4108",
      x"8748" & x"5595" & '0' & '0' & '1' & x"4343",
      x"2956" & x"3640" & '0' & '0' & '0' & x"6596",
      x"3414" & x"8526" & '1' & '0' & '1' & x"1941",
      x"4675" & x"7744" & '1' & '0' & '1' & x"2420",
      x"0200" & x"2955" & '1' & '0' & '0' & x"3156",
      x"9598" & x"4929" & '1' & '1' & '0' & x"4668",
      x"0425" & x"3750" & '1' & '1' & '1' & x"6674",
      x"7476" & x"7797" & '1' & '0' & '1' & x"5274",
      x"8599" & x"0241" & '0' & '1' & '0' & x"8358",
      x"0895" & x"0852" & '1' & '1' & '0' & x"0042",
      x"8380" & x"9204" & '0' & '0' & '1' & x"7584",
      x"6418" & x"5694" & '1' & '0' & '1' & x"2113",
      x"4091" & x"2375" & '1' & '1' & '0' & x"1715",
      x"5932" & x"3341" & '0' & '1' & '0' & x"2591",
      x"9240" & x"6179" & '0' & '0' & '1' & x"5419",
      x"0276" & x"4312" & '0' & '0' & '0' & x"4588",
      x"8623" & x"4084" & '0' & '0' & '1' & x"2707",
      x"9595" & x"8086" & '0' & '1' & '0' & x"1509",
      x"3966" & x"1513" & '1' & '0' & '0' & x"5480",
      x"5940" & x"1382" & '1' & '0' & '0' & x"7323",
      x"5050" & x"2039" & '1' & '1' & '0' & x"3010",
      x"7149" & x"6915" & '1' & '1' & '0' & x"0233",
      x"7791" & x"3660" & '1' & '0' & '1' & x"1452",
      x"2128" & x"1513" & '1' & '1' & '0' & x"0614",
      x"0096" & x"5652" & '1' & '0' & '0' & x"5749",
      x"4747" & x"7006" & '0' & '1' & '1' & x"7741",
      x"3744" & x"4135" & '0' & '1' & '1' & x"9609",
      x"8364" & x"8915" & '0' & '1' & '1' & x"9449",
      x"0763" & x"3697" & '1' & '0' & '0' & x"4461",
      x"6804" & x"1795" & '0' & '1' & '0' & x"5009",
      x"2316" & x"3616" & '1' & '0' & '0' & x"5933",
      x"0289" & x"2178" & '0' & '1' & '1' & x"8111",
      x"4226" & x"5342" & '0' & '0' & '0' & x"9568",
      x"2121" & x"7227" & '1' & '0' & '0' & x"9349",
      x"2285" & x"5633" & '1' & '0' & '0' & x"7919",
      x"8695" & x"2670" & '0' & '1' & '0' & x"6025",
      x"3149" & x"6169" & '0' & '1' & '1' & x"6980",
      x"3350" & x"0564" & '1' & '1' & '0' & x"2785",
      x"4344" & x"3383" & '1' & '1' & '0' & x"0960",
      x"0479" & x"0912" & '1' & '0' & '0' & x"1392",
      x"0048" & x"5988" & '1' & '1' & '1' & x"4059",
      x"3301" & x"5798" & '1' & '1' & '1' & x"7502",
      x"7520" & x"5415" & '1' & '1' & '0' & x"2104",
      x"7274" & x"4303" & '1' & '1' & '0' & x"2970",
      x"7765" & x"0204" & '1' & '1' & '0' & x"7560",
      x"5535" & x"5173" & '0' & '1' & '0' & x"0362",
      x"2087" & x"2976" & '0' & '1' & '1' & x"9111",
      x"5125" & x"9299" & '0' & '1' & '1' & x"5826",
      x"0979" & x"7725" & '1' & '0' & '0' & x"8705",
      x"8089" & x"4469" & '0' & '0' & '1' & x"2558",
      x"8949" & x"9025" & '1' & '1' & '1' & x"9923",
      x"9957" & x"7738" & '0' & '0' & '1' & x"7695",
      x"0185" & x"9827" & '0' & '1' & '1' & x"0358",
      x"2889" & x"6311" & '1' & '0' & '0' & x"9201",
      x"7769" & x"8540" & '0' & '1' & '1' & x"9229",
      x"1328" & x"3500" & '0' & '0' & '0' & x"4828",
      x"3845" & x"3059" & '0' & '0' & '0' & x"6904",
      x"5116" & x"2627" & '0' & '0' & '0' & x"7743",
      x"8612" & x"6188" & '0' & '0' & '1' & x"4800",
      x"9561" & x"6584" & '0' & '1' & '0' & x"2977",
      x"9087" & x"7036" & '0' & '0' & '1' & x"6123",
      x"6402" & x"5902" & '1' & '1' & '0' & x"0499",
      x"0276" & x"5416" & '0' & '1' & '1' & x"4860",
      x"4173" & x"8018" & '1' & '1' & '1' & x"6154",
      x"7241" & x"8305" & '0' & '0' & '1' & x"5546",
      x"5724" & x"1025" & '1' & '1' & '0' & x"4698",
      x"9411" & x"8565" & '0' & '0' & '1' & x"7976",
      x"7624" & x"8503" & '0' & '0' & '1' & x"6127",
      x"2607" & x"3804" & '0' & '0' & '0' & x"6411",
      x"2698" & x"9281" & '0' & '0' & '1' & x"1979",
      x"9830" & x"2935" & '0' & '1' & '0' & x"6895",
      x"8005" & x"3809" & '0' & '1' & '0' & x"4196",
      x"2698" & x"2582" & '0' & '1' & '0' & x"0116",
      x"2169" & x"2946" & '1' & '0' & '0' & x"5116",
      x"9965" & x"7074" & '0' & '0' & '1' & x"7039",
      x"2588" & x"0183" & '0' & '1' & '0' & x"2405",
      x"2027" & x"9975" & '0' & '1' & '1' & x"2052",
      x"4838" & x"9221" & '1' & '0' & '1' & x"4060",
      x"3321" & x"4048" & '1' & '0' & '0' & x"7370",
      x"5129" & x"2643" & '1' & '1' & '0' & x"2485",
      x"7940" & x"2194" & '1' & '1' & '0' & x"5745",
      x"9199" & x"5875" & '0' & '1' & '0' & x"3324",
      x"9949" & x"7657" & '0' & '1' & '0' & x"2292",
      x"0185" & x"9694" & '1' & '1' & '1' & x"0490",
      x"4966" & x"4578" & '1' & '0' & '0' & x"9545",
      x"5481" & x"2964" & '1' & '1' & '0' & x"2516",
      x"1591" & x"8049" & '0' & '0' & '0' & x"9640",
      x"6138" & x"5300" & '1' & '0' & '1' & x"1439",
      x"8138" & x"9419" & '0' & '0' & '1' & x"7557",
      x"3060" & x"6763" & '0' & '1' & '1' & x"6297",
      x"2470" & x"2756" & '0' & '1' & '1' & x"9714",
      x"1692" & x"2186" & '0' & '1' & '1' & x"9506",
      x"7915" & x"5222" & '1' & '1' & '0' & x"2692",
      x"2828" & x"9138" & '0' & '1' & '1' & x"3690",
      x"4172" & x"5450" & '1' & '1' & '1' & x"8721",
      x"2152" & x"2804" & '0' & '1' & '1' & x"9348",
      x"8217" & x"1811" & '0' & '1' & '0' & x"6406",
      x"0923" & x"4333" & '1' & '0' & '0' & x"5257",
      x"5716" & x"7743" & '0' & '1' & '1' & x"7973",
      x"0650" & x"2791" & '0' & '0' & '0' & x"3441",
      x"4489" & x"9800" & '1' & '0' & '1' & x"4290",
      x"3648" & x"1617" & '0' & '1' & '0' & x"2031",
      x"3712" & x"9693" & '0' & '1' & '1' & x"4019",
      x"7475" & x"6835" & '0' & '0' & '1' & x"4310",
      x"9648" & x"2249" & '1' & '0' & '1' & x"1898"
   );
 
begin

   uut: BCD_AddSub generic map (4) port map (A, B, cbi, sub, cbo, sum);

   process
   begin
      for i in test_vector'Range loop
      
         -- Assign test inputs
         A <= test_vector(i)(50 downto 35);
         B <= test_vector(i)(34 downto 19);
         cbi <= test_vector(i)(18);
         sub <= test_vector(i)(17);
         
         -- Compare outputs to expected values
         wait for 2ns;
         assert (cbo = test_vector(i)(16) and sum = test_vector(i)(15 downto 0))
            report "***** Test failed. *****"
            severity Failure;
      end loop;
      
      -- All tests are successful if we get this far
      report "***** All tests completed successfully. *****";
      wait;
   end process;

end testbench;
